package common is
    
    type queue_t is array(0 to 399) of integer range -300 to 600;
    
end package common;