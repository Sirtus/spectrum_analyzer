library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.common.all;
use work.trigonometric.all;

entity dft_test is
    port (
        clk: in std_logic;
        res: inout queue_t
    );
end entity dft_test; 

architecture arch of dft_test is
    -- constant data: queue_t := (
    --     0 , 7 , 13 , 19 , 25 , 31 , 37 , 43 , 48 , 54 , 59 , 64 , 69 , 73 , 77 , 81 ,           
    -- 85 , 88 , 91 , 93 , 95 , 97 , 99 , 100 , 100 , 100 , 100 , 100 , 99 , 98 , 96 , 94 , 91 , 89 ,
    --  86 , 82 , 78 , 74 , 70 , 65 , 60 , 55 , 50 , 44 , 39 , 33 , 27 , 21 , 15 , 8 , 2 , -4 , -10 , 
    --  -17 , -23 , -29 , -35 , -40 , -46 , -51 , -57 , -62 , -66 , -71 , -75 , -79 , -83 , -86 , -89 , 
    --  -92 , -94 , -96 , -97 , -98 , -99 , -99 , -99 , -99 , -98 , -97 , -95 , -93 , -91 , -88 , -85 ,
    --  -82 , -78 , -74 , -70 , -65 , -61 , -56 , -50 , -45 , -39 , -33 , -27 , -21 , -15 , -9 , -3 , 3 ,
    --   10 , 16 , 22 , 28 , 34 , 40 , 46 , 51 , 56 , 61 , 66 , 71 , 75 , 79 , 83 , 86 , 89 , 92 , 94 , 
    --   96 , 98 , 99 , 100 , 100 , 100 , 100 , 99 , 98 , 97 , 95 , 93 , 90 , 87 , 84 , 80 , 76 , 72 , 68 ,
    --   63 , 58 , 53 , 47 , 42 , 36 , 30 , 24 , 18 , 12 , 5 , -1 , -7 , -13 , -19 , -25 , -31 , -37 , -43 ,
    --   -49 , -54 , -59 , -64 , -69 , -73 , -77 , -81 , -84 , -87 , -90 , -93 , -95 , -96 , -98 , -99 , -99 ,
    --    -99 , -99 , -99 , -98 , -96 , -95 , -92 , -90 , -87 , -84 , -80 , -77 , -72 , -68 , -63 , -58 , -53 , 
    --    -48 , -42 , -36 , -31 , -25 , -19 , -12 , -6 , 0 , 6 , 13 , 19 , 25 , 31 , 37 , 43 , 48 , 54 , 59 , 64 ,
    --     68 , 73 , 77 , 81 , 84 , 88 , 91 , 93 , 95 , 97 , 99 , 100 , 100 , 100 , 100 , 100 , 99 , 98 , 96 , 94 , 
    --     92 , 89 , 86 , 82 , 79 , 74 , 70 , 66 , 61 , 56 , 50 , 45 , 39 , 33 , 27 , 21 , 15 , 9 , 3 , -4 , -10 , -16 , 
    --     -22, others => 0 );

    constant data: queue_t := (
        0, 10, 19, 27, 35, 42, 48, 53, 57, 60, 62, 62, 62, 61, 59, 57, 55, 53, 51, 49, 48, 46, 46, 46, 46, 46, 47, 48, 49, 50, 51, 52, 52, 52, 52, 51, 50, 49, 
        47, 46, 44, 43, 41, 40, 39, 38, 37, 36, 35, 34, 33, 32, 30, 27, 24, 20, 15, 9, 3, -4, -11, -19, -27, -34, -42, -49, -55, -61, -65, -68, -70, -71, -70, 
        -69, -66, -62, -57, -52, -47, -42, -36, -31, -27, -23, -20, -17, -16, -15, -15, -15, -16, -17, -18, -20, -21, -21, -22, -22, -21, -19, -18, -15, -12, -9,
         -6, -2, 1, 5, 9, 12, 15, 18, 21, 24, 27, 30, 33, 36, 40, 43, 47, 51, 56, 60, 65, 69, 73, 77, 80, 83, 85, 86, 85, 84, 81, 78, 73, 68, 62, 55, 48, 41, 34, 
        28, 21, 16, 12, 8, 6, 4, 4, 4, 5, 7, 9, 11, 13, 15, 17, 18, 18, 18, 17, 15, 12, 9, 5, 1, -4, -9, -14, -18, -23, -27, -31, -34, -36, -38, -40, -41, -42, 
        -43, -44, -44, -44, -44, -44, -45, -44, -44, -44, -43, -42, -40, -38, -35, -32, -28, -23, -17, -11, -5, 2, 8, 15, 21, 26, 31, 35, 39, 41, 42, 42, 41, 39,
         37, 33, 30, 26, 23, 19, 16, 14, 13, 12, 12, 14, 16, 19, 22, 26, 31, 35, 39, 44, 47, 51, 53, 55, 55, 55, 54, 52, 50, 47, 43, 39, 35, 31, 27, 23, 19, 15, 
        11, 7, 4, 0, -3, -6, -10, -14, -18, -22, -26, -30, -34, -38, -42, -46, -49, -51, -53, -54, -54, -54, -52, -50, -46, -43, -38, -34, -30, -25, -21, -18, 
        -15, -13, -11, -11, -12, -13, -15, -18, -22, -25, -29, -32, -36, -38, -40, -41, -41, -40, -38, -34, -30, -25, -20, -14, -7, -1, 6, 12, 18, 24, 29, 33, 
        36, 39, 41, 43, 44, 45, 45, 45, 46, 45, 45, 45, 45, 45, 44, 43, 42, 41, 39, 37, 35, 32, 28, 24, 19, 15, 10, 5, 0, -4, -8, -11, -14, -16, -17, -17, -17, 
        -16, -14, -12, -10, -8, -6, -4, -3, -3, -3, -5, -7, -11, -15, -20, -27, -33, -40, -47, -54, -61, -67, -72, -77, -80, -83, -84, -85, -84, -82, -80, -76, 
        -72, -68, -64, -59, -55, -50, -46, -42, -39, -35, -32, -29, -26, -23, -20, -17, -14, -11, -8, -4, 0, 3, 7, 10, 13, 16, 19, 20, 22, 23, 23, 22, 22, 21, 
        19, 18, 17, 16, 16, 16, 17, 18, 21, 24, 28, 32, 37, 43, 48, 53, 58, 63, 67, 70, 71, 72, 71, 69, 66, 62, 56, 50, 43, 35, 28, 20, 12, 5, -2, -8, -14, -19, 
        -23, -26, -29, -31, -32, -33, -34, -35, -36, -37, -38, -39, -40, -42, -43, -45, -46, -48, -49, -50, -51, -51, -51, -51, -50, -49, -48, -47, -46, -45, 
        -45, -45, -45, -45, -47, -48, -50, -52, -54, -56, -58, -60, -61, -61, -61, -59, -56, -52, -47, -41, -34, -26, -18, -9, others => 0
    );
    
    signal rout: queue_t := (others => 0);
begin

    p : process(clk)
    variable q: queue_t := (others => 0);
    begin
        if rising_edge(clk) then
            q := (others => 0);

            for i in 0 to 512 loop
                for j in 0 to 512 loop
                    q(i) := q(i) + (data(j) * app_sin((628*i*j)/5120));
                    
                end loop;
                rout(i) <= 300 - q(i)/3000;
            end loop;  
            -- rout <= q;

            
        end if;
        
    end process;
    
    -- g: for i in 0 to 10 generate
    --     gf: for j in 0 to 10 generate
    --         rout(i*10 + j) <= j when j < 600 else 600 - j;
    --     end generate gf;
    -- end generate g;
    res <= rout;
end architecture arch;