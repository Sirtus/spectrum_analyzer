package trigonometric is

    function apprrox_sin(x: integer) return integer;;
    
end package;

package body trigonometric is
    function apprrox_sin(x: integer) return integer is
        begin
            
        end function
end package body;