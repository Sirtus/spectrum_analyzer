library IEEE;
library work;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.common.all;

entity spectrum_analyzer is
    port(
        clk: in std_logic;

        red, green, blue: out std_logic_vector(3 downto 0);
        h_sync, v_sync: out std_logic;
		  
		mic_vcc: out std_logic := '1';
		mic_gnd: out std_logic := '0';

        sel: out std_logic := '0';
        lrcl: out std_logic;
        din: in std_logic;
        sclk: out std_logic;
        switch: in std_logic
    );
end spectrum_analyzer;

architecture arch of spectrum_analyzer is

    signal video_on: std_logic := '0';
    signal pixel_x, pixel_y: integer range 0 to 2047 := 0;
    signal mclk: std_logic := '0';
    signal dd, l_data, r_data : std_logic_vector(23 downto 0);
    signal do, do_i: isignal_t := (others => 0);
    signal do_cos, do_next: osignal_t := (others => 0);
    signal wr_en, do_fft: std_logic := '1';
    signal do_i_cnt: integer := 0;
    signal data_pixel: std_logic_vector(15 downto 0) := (others => '0');
    signal data_pixel_int: integer := 0;
    
    signal done_f: std_logic := '0';
    signal ws: std_logic := '0';

    signal addressA, addressB: std_logic_vector(14 downto 0);
    signal dataA, dataB, qA, qB: std_logic_vector(15 downto 0);
    signal wrA, wrB: std_logic;
    
    signal last_column: integer;
    

    begin 

    bclk: entity work.bclk
    port map( inclk0 => clk, c0 => mclk);

    reg: entity work.shift_reg
    port map(clock => clk, address_a => addressA, address_b => addressB, data_a => dataA, 
             data_b => dataB, wren_a => wrA, wren_b => wrB, q_a => qA, q_b => qB);

    vga: entity work.vga_controller
    port map( clk => clk, video_on => video_on, pixel_x => pixel_x, pixel_y => pixel_y,
              h_sync => h_sync, v_sync => v_sync);

    plot: entity work.plot_controller
    port map(clk => clk, video_on => video_on, pixel_x => pixel_x, pixel_y => pixel_y, 
             red => red, green => green, blue => blue, do => data_pixel, last_column => last_column, addressA => addressA, qA => qA);

    
    fft: entity work.fft
    port map(clk => clk,  do_fft => switch, done => done_f, wr_en => wr_en, data_in => l_data, last_column => last_column, general_ram_addr => addressB, general_ram_data => dataB, general_ram_wren => wrB);


    -- process(clk)
    -- variable pixel_addr: unsigned(13 downto 0) := (others => '0'); 
    -- variable current_column: integer range 0 to 127 := 0;
    -- variable col_x, row_y: integer range 0 to 127 := 0;
    -- begin
    --     if rising_edge(clk) then
    --         if pixel_y <= 512 and pixel_x <= 128 then
    --             if pixel_x = 0 and pixel_y mod 8 = 0 then
    --                 row_y := row_y + 1;
    --             end if;
    --             col_y <= (current_column * N_DIV_2) + row_y;
    --             pixel_addr := to_unsigned(col_y, addressA'length);
    --             current_column := (last_column + col_x);
    --             addressA <= std_logic_vector(pixel_addr);
    --             data_pixel <= qA;
    --             if pixel_x mod 4 = 0 then
    --                 col_x := col_x + 1;
    --             end if;
    --         else
    --             col_x := 0;
    --             data_pixel <= (others => '0');
    --             if pixel_y >= 512 then
    --                 row_y := 0;
    --             end if;
    --         end if;
    --     end if;
    -- end process;

    -- do_fft <= '1'; --switch;

    i2s: entity work.i2s_receiver
    port map(sclk => mclk, ws => ws, d_rx => din, l_data => l_data, r_data => r_data, sel => sel,
    read_en => wr_en);

    lrcl <= ws;
    sclk <= mclk;
    wrA <= '0';
    dataA <= (others => '0');

end arch;

