package common is
    
    type queue_t is array(0 to 799) of integer range 0 to 600;
    
end package common;