library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.common.all;


entity fft_tb is
end fft_tb;

architecture sim of fft_tb is

    constant clk_period : time := 10 ps;

    signal clk : std_logic := '1';
    signal rst : std_logic := '1';

    signal res: queue_t := (others => 0);
    -- signal data: queue_t := 
    -- (
    --     0 , 9 , 19 , 29 , 38 , 47 , 56 , 64 , 71 , 78 , 
    --     84 , 89 , 93 , 96 , 98 , 99 , 99 , 99 , 97 , 94 , 
    --     90 , 86 , 80 , 74 , 67 , 59 , 51 , 42 , 33 , 23 , 
    --     14 , 4 
    -- );
    signal data: queue_t := 
    (
        -- 35, 35, 64, 106, 35, -106, -135, others => -35 
        -- 0, -106,  200 ,-106, 0 , 106, -200 , 106
        -- 170, 170, 199, 241, 170, 29, 0, 100
        -- 255,12, 123, 255, 3, 12, 255, 12
        -- 0, 1, 2, 3, 4, 5, 6, 7
        -- 0, -8, -154, 109, 161, 153, 171, -35, -122, -142, -147, -41, 198, 26, 57, 113, 
        -- -191, -168, 3, 136, 75, 178, -123, -163, 8, 193, 132, -117, -181, -139, -188, 
        -- 47, 1, -136, 193, 166, -20, -61, 119, -71, -197, -163, -186, -199, -189, -52, 
        -- 152, 146, -167, -8, 13, -125, 117, -126, 78, 181, 167, 131, -166, -185, -133, 
        -- -87, -145, -144, 182, 197, 42, -181, -133, -53, 112, -77, 167, 23, -138, -53, 
        -- 117, 197, 141, -84, -167, -28, 190, 186, -189, 193, 99, 182, -197, -96, -189, 
        -- -105, -20, -109, -189, -185, 0, 199, 192, 73, -181, -47, -183, 198, 8, 182, 
        -- -3, -136, 75, 162, -73, -185, -191, -175, -180, 111, 198, 41, -182, -86, -122, 
        -- 96, -197, -146, 161, 191, 200, 118, 1, -117, -199, -190, -160, 147, 198, -95, 
        -- 123, 87, 183, -40, -197, -110, 181, 176, 192, 186, 74, -161, -74, 137, 4, 
        -- -181, -7, -197, 184, 48, 182, -72, -191, -198, 0, 186, 190, 110, 21, 106, 
        -- 190, 97, 198, -181, -98, -192, 190, -185, -189, 29, 168, 85, -140, -196, -116, 
        -- 54, 139, -22, -166, 78, -111, 54, 134, 182, -41, -196, -181, 145, 146, 88, 
        -- 134, 186, 167, -130, -166, -180, -77, 127, -116, 126, -12, 9, 168, -145, -151, 
        -- 53, 190, 200, 187, 164, 198, 72, -118, 62, 21, -165, -192, 137, 1, -46, 
        -- 189, 140, 182, 118, -131, -192, -7, 164, 124, -177, -74, -135, -2, 169, 192, 
        -- -112, -56, -25, -197, 42, 148, 143, 123, 36, -170, -152, -160, -108, 155, 9, 
        0, -122, -191, 8, 1, -197, -167, 167, 182, 167, -167, -197, 0, 8, -191, -122, 
        1, 123, 192, -7, 0, 198, 168, -166, -181, -166, 168, 198, 1, -7, 192, 123, others => 0
    );
    -- signal do_next: queue_t := (others => 0);
    signal do_fft: std_logic := '1';
    signal done: std_logic := '0';

begin

    clk <= not clk after clk_period / 2;

    fft: entity work.fft
    port map(
        clk => clk,
        data_i => data,
        do_fft=> do_fft,
        done=> done,
        res=> res
    );


end architecture;