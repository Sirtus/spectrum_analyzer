module fft_top;
  import uvm_pkg::*;



  initial begin

  end
endmodule
