package common is
    
    type queue_t is array(0 to 255) of integer range -60000 to 60000;
--     type vec_t is array(0 to 799) of integer range 0 to 100;
	 
	 constant ccc: queue_t := (0 , 7 , 13 , 19 , 25 , 31 , 37 , 43 , 48 , 54 , 59 , 64 , 69 , 73 , 77 , 81 , 
     85 , 88 , 91 , 93 , 95 , 97 , 99 , 100 , 100 , 100 , 100 , 100 , 99 , 98 , 96 , 94 , 91 , 89 , 86 , 82 , 
     78 , 74 , 70 , 65 , 60 , 55 , 50 , 44 , 39 , 33 , 27 , 21 , 15 , 8 , 2 , -4 , -10 , -17 , -23 , -29 , -35 , 
     -40 , -46 , -51 , -57 , -62 , -66 , -71 , -75 , -79 , -83 , -86 , -89 , -92 , -94 , -96 , -97 , -98 , -99 , -99 , 
     -99 , -99 , -98 , -97 , -95 , -93 , -91 , -88 , -85 , -82 , -78 , -74 , -70 , -65 , -61 , -56 , -50 , -45 , -39 , 
     -33 , -27 , -21 , -15 , -9 , -3 , 3 , 10 , 16 , 22 , 28 , 34 , 40 , 46 , 51 , 56 , 61 , 66 , 71 , 75 , 79 , 83 , 86 , 
     89 , 92 , 94 , 96 , 98 , 99 , 100 , 100 , 100 , 100 , 99 , 98 , 97 , 95 , 93 , 90 , 87 , 84 , 80 , 76 , 72 , 68 , 63 , 
     58 , 53 , 47 , 42 , 36 , 30 , 24 , 18 , 12 , 5 , -1 , -7 , -13 , -19 , -25 , -31 , -37 , -43 , -49 , -54 , -59 , -64 , 
     -69 , -73 , -77 , -81 , -84 , -87 , -90 , -93 , -95 , -96 , -98 , -99 , -99 , -99 , -99 , -99 , -98 , -96 , -95 , -92 , 
     -90 , -87 , -84 , -80 , -77 , -72 , -68 , -63 , -58 , -53 , -48 , -42 , -36 , -31 , -25 , -19 , -12 , -6 , 0 , 6 , 13 , 
     19 , 25 , 31 , 37 , 43 , 48 , 54 , 59 , 64 , 68 , 73 , 77 , 81 , 84 , 88 , 91 , 93 , 95 , 97 , 99 , 100 , 100 , 100 , 100 , 
     100 , 99 , 98 , 96 , 94 , 92 , 89 , 86 , 82 , 79 , 74 , 70 , 66 , 61 , 56 , 50 , 45 , 39 , 33 , 27 , 21 , 15 , 9 , 3 , -4 , -10 , -16 , -22 );
     
-- 	(

--               0 , 13 , 26 , 38 , 50 , 61 , 72 , 81 , 89 , 96 , 101 , 105 , 107 , 107 , 107 , 104 , 
--               100 , 95 , 88 , 80 , 71 , 61 , 50 , 39 , 27 , 15 , 3 , -7 , -19 , -30 , -40 , -49 , 
--               -57 , -63 , -69 , -73 , -75 , -76 , -76 , -73 , -70 , -65 , -58 , -50 , -41 , -30 , -19 , -7 , 
--               4 , 17 , 30 , 44 , 56 , 69 , 81 , 92 , 102 , 112 , 120 , 126 , 131 , 135 , 137 , 138 , 
--               137 , 134 , 130 , 125 , 118 , 110 , 101 , 91 , 80 , 69 , 57 , 45 , 33 , 21 , 10 , 0 , 
--               -10 , -19 , -27 , -34 , -40 , -44 , -46 , -47 , -47 , -45 , -41 , -36 , -29 , -21 , -12 , -2 , 
--               8 , 20 , 32 , 45 , 58 , 71 , 84 , 97 , 108 , 120 , 130 , 139 , 147 , 153 , 158 , 162 , 
--               164 , 164 , 163 , 161 , 157 , 151 , 144 , 136 , 127 , 117 , 106 , 94 , 82 , 70 , 58 , 46 , 
--               35 , 24 , 14 , 4 , -3 , -10 , -15 , -20 , -22 , -23 , -23 , -21 , -18 , -13 , -6 , 1 , 
--               10 , 20 , 31 , 42 , 55 , 67 , 80 , 93 , 106 , 118 , 130 , 141 , 151 , 160 , 168 , 174 , 
--               179 , 182 , 184 , 185 , 183 , 181 , 176 , 171 , 164 , 155 , 146 , 136 , 125 , 113 , 101 , 89 , 
--               76 , 64 , 53 , 42 , 31 , 22 , 13 , 6 , 1 , -3 , -6 , -7 , -7 , -5 , -2 , 2 , 
--               9 , 16 , 25 , 35 , 46 , 57 , 69 , 82 , 95 , 107 , 120 , 132 , 144 , 154 , 164 , 173 , 
--               180 , 187 , 191 , 195 , 196 , 197 , 195 , 192 , 188 , 182 , 175 , 166 , 157 , 146 , 135 , 123 , 
--               111 , 98 , 86 , 74 , 62 , 50 , 40 , 30 , 22 , 14 , 9 , 4 , 1 , 0 , 0 , 1 , 
--               4 , 9 , 15 , 22 , 31 , 41 , 51 , 63 , 75 , 87 , 99 , 112 , 124 , 136 , 148 , 158

-- --        0 , 13 , 26 , 38 , 50 , 61 , 72 , 81 , 89 , 96 , 101 , 105 , 107 , 107 , 107 , 104 , 
-- -- 100 , 95 , 88 , 80 , 71 , 61 , 50 , 39 , 27 , 15 , 3 , -7 , -19 , -30 , -40 , -49 , 
-- -- -57 , -63 , -69 , -73 , -75 , -76 , -76 , -73 , -70 , -65 , -58 , -50 , -41 , -30 , -19 , -7 , 
-- -- 4 , 17 , 30 , 44 , 56 , 69 , 81 , 92 , 102 , 112 , 120 , 126 , 131 , 135 , 137 , 138 , 
-- -- 137 , 134 , 130 , 125 , 118 , 110 , 101 , 91 , 80 , 69 , 57 , 45 , 33 , 21 , 10 , 0 , 
-- -- -10 , -19 , -27 , -34 , -40 , -44 , -46 , -47 , -47 , -45 , -41 , -36 , -29 , -21 , -12 , -2 , 
-- -- 8 , 20 , 32 , 45 , 58 , 71 , 84 , 97 , 108 , 120 , 130 , 139 , 147 , 153 , 158 , 162 , 
-- -- 164 , 164 , 163 , 161 , 157 , 151 , 144 , 136 , 127 , 117 , 106 , 94 , 82 , 70 , 58 , 46 , 
-- -- 35 , 24 , 14 , 4 , -3 , -10 , -15 , -20 , -22 , -23 , -23 , -21 , -18 , -13 , -6 , 1 , 
-- -- 10 , 20 , 31 , 42 , 55 , 67 , 80 , 93 , 106 , 118 , 130 , 141 , 151 , 160 , 168 , 174 , 
-- -- 179 , 182 , 184 , 185 , 183 , 181 , 176 , 171 , 164 , 155 , 146 , 136 , 125 , 113 , 101 , 89 , 
-- -- 76 , 64 , 53 , 42 , 31 , 22 , 13 , 6 , 1 , -3 , -6 , -7 , -7 , -5 , -2 , 2 , 
-- -- 9 , 16 , 25 , 35 , 46 , 57 , 69 , 82 , 95 , 107 , 120 , 132 , 144 , 154 , 164 , 173 , 
-- -- 180 , 187 , 191 , 195 , 196 , 197 , 195 , 192 , 188 , 182 , 175 , 166 , 157 , 146 , 135 , 123 , 
-- -- 111 , 98 , 86 , 74 , 62 , 50 , 40 , 30 , 22 , 14 , 9 , 4 , 1 , 0 , 0 , 1 , 
-- -- 4 , 9 , 15 , 22 , 31 , 41 , 51 , 63 , 75 , 87 , 99 , 112 , 124 , 136 , 148 , 158 , 
-- -- 168 , 176 , 184 , 190 , 194 , 197 , 199 , 199 , 197 , 194 , 189 , 183 , 176 , 167 , 157 , 147 , 
-- -- 135 , 123 , 111 , 98 , 86 , 73 , 61 , 50 , 39 , 29 , 20 , 13 , 7 , 2 , 0 , -2 , 
-- -- -2 , -1 , 1 , 6 , 12 , 19 , 27 , 37 , 47 , 58 , 70 , 82 , 95 , 107 , 119 , 131 , 
-- -- 142 , 152 , 162 , 170 , 177 , 183 , 188 , 190 , 192 , 192 , 190 , 186 , 182 , 175 , 168 , 159 , 
-- -- 149 , 138 , 126 , 114 , 101 , 89 , 76 , 63 , 51 , 39 , 28 , 18 , 9 , 2 , -4 , -9 , 
-- -- -12 , -14 , -14 , -13 , -10 , -6 , 0 , 6 , 14 , 23 , 34 , 45 , 56 , 68 , 80 , 93 , 
-- -- 105 , 116 , 127 , 137 , 147 , 155 , 162 , 167 , 172 , 174 , 176 , 175 , 173 , 170 , 165 , 158 , 
-- -- 150 , 141 , 131 , 120 , 108 , 96 , 83 , 70 , 57 , 44 , 32 , 20 , 9 , 0 , -9 , -17 , 
-- -- -23 , -28 , -32 , -34 , -35 , -34 , -31 , -27 , -21 , -14 , -6 , 2 , 12 , 23 , 34 , 46 , 
-- -- 58 , 70 , 82 , 94 , 104 , 114 , 124 , 132 , 139 , 144 , 148 , 151 , 152 , 151 , 149 , 146 , 
-- -- 140 , 134 , 126 , 117 , 106 , 95 , 83 , 71 , 58 , 45 , 32 , 19 , 6 , -5 , -16 , -26 , 
-- -- -35 , -43 , -50 , -55 , -59 , -61 , -61 , -60 , -58 , -54 , -48 , -41 , -33 , -24 , -14 , -4 , 
-- -- 7 , 18 , 30 , 42 , 54 , 65 , 76 , 86 , 95 , 103 , 110 , 115 , 119 , 122 , 123 , 122 , 
-- -- 120 , 116 , 111 , 105 , 97 , 87 , 77 , 66 , 54 , 41 , 28 , 15 , 2 , -10 , -23 , -35 , 
-- -- -46 , -56 , -65 , -73 , -80 , -85 , -89 , -91 , -92 , -91 , -88 , -84 , -79 , -72 , -64 , -55 , 
-- -- -45 , -34 , -23 , -11 , 0 , 11 , 23 , 34 , 45 , 55 , 64 , 72 , 79 , 84 , 88 , 91 , 
-- -- 92 , 91 , 89 , 85 , 80 , 73 , 65 , 56 , 46 , 35 , 23 , 10 , -2 , -15 , -28 , -41 , 
-- -- -54 , -66 , -77 , -87 , -97 , -105 , -111 , -116 , -120 , -122 , -123 , -122 , -119 , -115 , -110 , -103 , 
-- -- -95 , -86 , -76 , -65 , -54 , -42 , -30 , -18 , -7 , 4 , 14 , 24 , 33 , 41 , 48 , 54 , 
-- -- 58 , 60 , 61 , 61 , 59 , 55 , 50 , 43 , 35 , 26 , 16 , 5 , -6 , -19 , -32 , -45 , 
-- -- -58 , -71 , -83 , -95 , -106 , -117 , -126 , -134 , -140 , -146 , -149 , -151 , -152 , -151 , -148 , -144 , 
-- -- -139 , -132 , -124 , -114 , -104 , -94 , -82 , -70 , -58 , -46 , -34 , -23 , -12 , -2 , 6 , 14 , 
-- -- 21 , 27 , 31 , 34 , 35 , 34 , 32 , 28 , 23 , 17 , 9 , 0 , -9 , -20 , -32 , -44 , 
-- -- -57 , -70 , -83 , -96 , -108 , -120 , -131 , -141 , -150 , -158 , -165 , -170 , -173 , -175 , -176 , -174 , 
-- -- -172 , -167 , -162 , -155 , -147 , -137 , -127 , -116 , -105 , -93 , -80 , -68 , -56 , -45 , -34 , -23 , 
-- -- -14 , -6 , 0 , 6 , 10 , 13 , 14 , 14 , 12 , 9 , 4 , -2 , -9 , -18 , -28 , -39 , 
-- -- -51 , -63 , -76 , -89 , -101 , -114 , -126 , -138 , -149 , -159 , -168 , -175 , -182 , -186 , -190 , -192 , 
-- -- -192 , -190 , -188 , -183 , -177 , -170 , -162 , -152 , -142 , -131 , -119 , -107 , -95 , -82 , -70 , -58 , 
-- -- -47 , -37 , -27 , -19 , -12 , -6 , -1 , 1 , 2 , 2 , 0 , -2 , -7 , -13 , -20 , -29 , 
-- -- -39 , -50 , -61 , -73 , -86 , -98 , -111 , -123 , -135 , -147 , -157 , -167 , -176 , -183 , -189 , -194 , 
-- -- -197 , -199 , -199 , -197 , -194 , -190 , -184 , -176 , -168 , -158 , -148 , -136 , -124 , -112 , -100 , -87 , 
-- -- -75 , -63 , -51 , -41 , -31 , -22 , -15 , -9 , -4 , -1 , 0 , 0 , -1 , -4 , -9 , -14 , 
-- -- -22 , -30 , -40 , -50 , -62 , -74 , -86 , -98 , -111 , -123 , -135 , -146 , -157 , -166 , -175 , -182 , 
-- -- -188 , -192 , -195 , -197 , -196 , -195 , -191 , -187 , -180 , -173 , -164 , -154 , -144 , -132 , -120 , -107
-- 	); 
    
end package common;