package i2s_pkg;
    `include "../tests/i2s_test.svh"
endpackage
