package common is
    
    type queue_t is array(0 to 799) of integer;
    
end package common;